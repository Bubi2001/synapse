module ALU (
    input  logic        clk,
    input  logic        rst_n,
    input  logic [6:0]  opcode,
    input  logic [31:0] opA,
    input  logic [31:0] opB,
    input  logic        cin,
    input  logic        busEnable,
    output logic [31:0] aluOut,
    output logic [4:0]  flags
)



endmodule