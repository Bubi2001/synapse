package FPUOperations;
    // Define an enum for FPU operations
    typedef enum logic [5:0] {
        FPU_NOP         = 6'h00,
        FPU_ADD_S       = 6'h01,
        FPU_SUB_S       = 6'h02,
        FPU_MUL_S       = 6'h03,
        FPU_DIV_S       = 6'h04,
        FPU_MIN_S       = 6'h05,
        FPU_MAX_S       = 6'h06,
        FPU_SQRT_S      = 6'h07,
        FPU_MADD_S      = 6'h08,
        FPU_MSUB_S      = 6'h09,
        FPU_NMADD_S     = 6'h0A,
        FPU_NMSUB_S     = 6'h0B,
        FPU_CVT_W_S     = 6'h0C,
        FPU_CVT_WU_S    = 6'h0D,
        FPU_CVT_S_W     = 6'h0E,
        FPU_CVT_S_WU    = 6'h0F,
        FPU_SGNJ_S      = 6'h10,
        FPU_SGNJN_S     = 6'h11,
        FPU_SGNJX_S     = 6'h12,
        FPU_EQ_S        = 6'h13,
        FPU_LT_S        = 6'h14,
        FPU_LE_S        = 6'h15,
        FPU_ADD_D       = 6'h16,
        FPU_SUB_D       = 6'h17,
        FPU_MUL_D       = 6'h18,
        FPU_DIV_D       = 6'h19,
        FPU_MIN_D       = 6'h1A,
        FPU_MAX_D       = 6'h1B,
        FPU_SQRT_D      = 6'h1C,
        FPU_MADD_D      = 6'h1D,
        FPU_MSUB_D      = 6'h1E,
        FPU_NMADD_D     = 6'h1F,
        FPU_NMSUB_D     = 6'h20,
        FPU_CVT_S_D     = 6'h21,
        FPU_CVT_D_S     = 6'h22,
        FPU_CVT_W_D     = 6'h23,
        FPU_CVT_WU_D    = 6'h24,
        FPU_CVT_D_W     = 6'h25,
        FPU_CVT_D_WU    = 6'h26,
        FPU_SGNJ_D      = 6'h27,
        FPU_SGNJN_D     = 6'h28,
        FPU_SGNJX_D     = 6'h29,
        FPU_EQ_D        = 6'h2A,
        FPU_LT_D        = 6'h2B,
        FPU_LE_D        = 6'h2C
    } fpu_op_t;
endpackage
