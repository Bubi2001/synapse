module Synapse (
    input  logic        clk,
    input  logic        rst_n
);
    
endmodule